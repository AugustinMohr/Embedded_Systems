-- soc_system.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity soc_system is
	port (
		clk_clk                                     : in    std_logic                     := '0';             --                          clk.clk
		hps_0_ddr_mem_a                             : out   std_logic_vector(14 downto 0);                    --                    hps_0_ddr.mem_a
		hps_0_ddr_mem_ba                            : out   std_logic_vector(2 downto 0);                     --                             .mem_ba
		hps_0_ddr_mem_ck                            : out   std_logic;                                        --                             .mem_ck
		hps_0_ddr_mem_ck_n                          : out   std_logic;                                        --                             .mem_ck_n
		hps_0_ddr_mem_cke                           : out   std_logic;                                        --                             .mem_cke
		hps_0_ddr_mem_cs_n                          : out   std_logic;                                        --                             .mem_cs_n
		hps_0_ddr_mem_ras_n                         : out   std_logic;                                        --                             .mem_ras_n
		hps_0_ddr_mem_cas_n                         : out   std_logic;                                        --                             .mem_cas_n
		hps_0_ddr_mem_we_n                          : out   std_logic;                                        --                             .mem_we_n
		hps_0_ddr_mem_reset_n                       : out   std_logic;                                        --                             .mem_reset_n
		hps_0_ddr_mem_dq                            : inout std_logic_vector(31 downto 0) := (others => '0'); --                             .mem_dq
		hps_0_ddr_mem_dqs                           : inout std_logic_vector(3 downto 0)  := (others => '0'); --                             .mem_dqs
		hps_0_ddr_mem_dqs_n                         : inout std_logic_vector(3 downto 0)  := (others => '0'); --                             .mem_dqs_n
		hps_0_ddr_mem_odt                           : out   std_logic;                                        --                             .mem_odt
		hps_0_ddr_mem_dm                            : out   std_logic_vector(3 downto 0);                     --                             .mem_dm
		hps_0_ddr_oct_rzqin                         : in    std_logic                     := '0';             --                             .oct_rzqin
		hps_0_io_hps_io_emac1_inst_TX_CLK           : out   std_logic;                                        --                     hps_0_io.hps_io_emac1_inst_TX_CLK
		hps_0_io_hps_io_emac1_inst_TXD0             : out   std_logic;                                        --                             .hps_io_emac1_inst_TXD0
		hps_0_io_hps_io_emac1_inst_TXD1             : out   std_logic;                                        --                             .hps_io_emac1_inst_TXD1
		hps_0_io_hps_io_emac1_inst_TXD2             : out   std_logic;                                        --                             .hps_io_emac1_inst_TXD2
		hps_0_io_hps_io_emac1_inst_TXD3             : out   std_logic;                                        --                             .hps_io_emac1_inst_TXD3
		hps_0_io_hps_io_emac1_inst_RXD0             : in    std_logic                     := '0';             --                             .hps_io_emac1_inst_RXD0
		hps_0_io_hps_io_emac1_inst_MDIO             : inout std_logic                     := '0';             --                             .hps_io_emac1_inst_MDIO
		hps_0_io_hps_io_emac1_inst_MDC              : out   std_logic;                                        --                             .hps_io_emac1_inst_MDC
		hps_0_io_hps_io_emac1_inst_RX_CTL           : in    std_logic                     := '0';             --                             .hps_io_emac1_inst_RX_CTL
		hps_0_io_hps_io_emac1_inst_TX_CTL           : out   std_logic;                                        --                             .hps_io_emac1_inst_TX_CTL
		hps_0_io_hps_io_emac1_inst_RX_CLK           : in    std_logic                     := '0';             --                             .hps_io_emac1_inst_RX_CLK
		hps_0_io_hps_io_emac1_inst_RXD1             : in    std_logic                     := '0';             --                             .hps_io_emac1_inst_RXD1
		hps_0_io_hps_io_emac1_inst_RXD2             : in    std_logic                     := '0';             --                             .hps_io_emac1_inst_RXD2
		hps_0_io_hps_io_emac1_inst_RXD3             : in    std_logic                     := '0';             --                             .hps_io_emac1_inst_RXD3
		hps_0_io_hps_io_sdio_inst_CMD               : inout std_logic                     := '0';             --                             .hps_io_sdio_inst_CMD
		hps_0_io_hps_io_sdio_inst_D0                : inout std_logic                     := '0';             --                             .hps_io_sdio_inst_D0
		hps_0_io_hps_io_sdio_inst_D1                : inout std_logic                     := '0';             --                             .hps_io_sdio_inst_D1
		hps_0_io_hps_io_sdio_inst_CLK               : out   std_logic;                                        --                             .hps_io_sdio_inst_CLK
		hps_0_io_hps_io_sdio_inst_D2                : inout std_logic                     := '0';             --                             .hps_io_sdio_inst_D2
		hps_0_io_hps_io_sdio_inst_D3                : inout std_logic                     := '0';             --                             .hps_io_sdio_inst_D3
		hps_0_io_hps_io_usb1_inst_D0                : inout std_logic                     := '0';             --                             .hps_io_usb1_inst_D0
		hps_0_io_hps_io_usb1_inst_D1                : inout std_logic                     := '0';             --                             .hps_io_usb1_inst_D1
		hps_0_io_hps_io_usb1_inst_D2                : inout std_logic                     := '0';             --                             .hps_io_usb1_inst_D2
		hps_0_io_hps_io_usb1_inst_D3                : inout std_logic                     := '0';             --                             .hps_io_usb1_inst_D3
		hps_0_io_hps_io_usb1_inst_D4                : inout std_logic                     := '0';             --                             .hps_io_usb1_inst_D4
		hps_0_io_hps_io_usb1_inst_D5                : inout std_logic                     := '0';             --                             .hps_io_usb1_inst_D5
		hps_0_io_hps_io_usb1_inst_D6                : inout std_logic                     := '0';             --                             .hps_io_usb1_inst_D6
		hps_0_io_hps_io_usb1_inst_D7                : inout std_logic                     := '0';             --                             .hps_io_usb1_inst_D7
		hps_0_io_hps_io_usb1_inst_CLK               : in    std_logic                     := '0';             --                             .hps_io_usb1_inst_CLK
		hps_0_io_hps_io_usb1_inst_STP               : out   std_logic;                                        --                             .hps_io_usb1_inst_STP
		hps_0_io_hps_io_usb1_inst_DIR               : in    std_logic                     := '0';             --                             .hps_io_usb1_inst_DIR
		hps_0_io_hps_io_usb1_inst_NXT               : in    std_logic                     := '0';             --                             .hps_io_usb1_inst_NXT
		hps_0_io_hps_io_spim1_inst_CLK              : out   std_logic;                                        --                             .hps_io_spim1_inst_CLK
		hps_0_io_hps_io_spim1_inst_MOSI             : out   std_logic;                                        --                             .hps_io_spim1_inst_MOSI
		hps_0_io_hps_io_spim1_inst_MISO             : in    std_logic                     := '0';             --                             .hps_io_spim1_inst_MISO
		hps_0_io_hps_io_spim1_inst_SS0              : out   std_logic;                                        --                             .hps_io_spim1_inst_SS0
		hps_0_io_hps_io_uart0_inst_RX               : in    std_logic                     := '0';             --                             .hps_io_uart0_inst_RX
		hps_0_io_hps_io_uart0_inst_TX               : out   std_logic;                                        --                             .hps_io_uart0_inst_TX
		hps_0_io_hps_io_i2c0_inst_SDA               : inout std_logic                     := '0';             --                             .hps_io_i2c0_inst_SDA
		hps_0_io_hps_io_i2c0_inst_SCL               : inout std_logic                     := '0';             --                             .hps_io_i2c0_inst_SCL
		hps_0_io_hps_io_i2c1_inst_SDA               : inout std_logic                     := '0';             --                             .hps_io_i2c1_inst_SDA
		hps_0_io_hps_io_i2c1_inst_SCL               : inout std_logic                     := '0';             --                             .hps_io_i2c1_inst_SCL
		hps_0_io_hps_io_gpio_inst_GPIO09            : inout std_logic                     := '0';             --                             .hps_io_gpio_inst_GPIO09
		hps_0_io_hps_io_gpio_inst_GPIO35            : inout std_logic                     := '0';             --                             .hps_io_gpio_inst_GPIO35
		hps_0_io_hps_io_gpio_inst_GPIO40            : inout std_logic                     := '0';             --                             .hps_io_gpio_inst_GPIO40
		hps_0_io_hps_io_gpio_inst_GPIO53            : inout std_logic                     := '0';             --                             .hps_io_gpio_inst_GPIO53
		hps_0_io_hps_io_gpio_inst_GPIO54            : inout std_logic                     := '0';             --                             .hps_io_gpio_inst_GPIO54
		hps_0_io_hps_io_gpio_inst_GPIO61            : inout std_logic                     := '0';             --                             .hps_io_gpio_inst_GPIO61
		lcd_controller_0_conduit_end_export_cs_n    : out   std_logic;                                        -- lcd_controller_0_conduit_end.export_cs_n
		lcd_controller_0_conduit_end_export_data    : out   std_logic_vector(15 downto 0);                    --                             .export_data
		lcd_controller_0_conduit_end_export_d_c_n   : out   std_logic;                                        --                             .export_d_c_n
		lcd_controller_0_conduit_end_export_lcd_on  : out   std_logic;                                        --                             .export_lcd_on
		lcd_controller_0_conduit_end_export_rd_n    : out   std_logic;                                        --                             .export_rd_n
		lcd_controller_0_conduit_end_export_reset_n : out   std_logic;                                        --                             .export_reset_n
		lcd_controller_0_conduit_end_export_wr_n    : out   std_logic;                                        --                             .export_wr_n
		pio_leds_external_connection_export         : out   std_logic_vector(7 downto 0);                     -- pio_leds_external_connection.export
		reset_reset_n                               : in    std_logic                     := '0'              --                        reset.reset_n
	);
end entity soc_system;

architecture rtl of soc_system is
	component LT24_controller is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			nReset         : in  std_logic                     := 'X';             -- reset_n
			AM_address     : out std_logic_vector(31 downto 0);                    -- address
			AM_read        : out std_logic;                                        -- read
			AM_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			AM_waitRQ      : in  std_logic                     := 'X';             -- waitrequest
			AM_BurstCount  : out std_logic_vector(7 downto 0);                     -- burstcount
			AM_Rddatavalid : in  std_logic                     := 'X';             -- readdatavalid
			CS_N           : out std_logic;                                        -- export_cs_n
			DATA           : out std_logic_vector(15 downto 0);                    -- export_data
			D_C_N          : out std_logic;                                        -- export_d_c_n
			LCD_ON         : out std_logic;                                        -- export_lcd_on
			RD_N           : out std_logic;                                        -- export_rd_n
			RESET_N        : out std_logic;                                        -- export_reset_n
			WR_N           : out std_logic;                                        -- export_wr_n
			AS_address     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			AS_write       : in  std_logic                     := 'X';             -- write
			AS_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			AS_read        : in  std_logic                     := 'X';             -- read
			AS_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			AS_CS          : in  std_logic                     := 'X';             -- chipselect
			AS_irq         : out std_logic                                         -- irq
		);
	end component LT24_controller;

	component altera_address_span_extender is
		generic (
			DATA_WIDTH           : integer                       := 32;
			BYTEENABLE_WIDTH     : integer                       := 4;
			MASTER_ADDRESS_WIDTH : integer                       := 32;
			SLAVE_ADDRESS_WIDTH  : integer                       := 16;
			SLAVE_ADDRESS_SHIFT  : integer                       := 2;
			BURSTCOUNT_WIDTH     : integer                       := 1;
			CNTL_ADDRESS_WIDTH   : integer                       := 1;
			SUB_WINDOW_COUNT     : integer                       := 1;
			MASTER_ADDRESS_DEF   : std_logic_vector(63 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000"
		);
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			avs_s0_address       : in  std_logic_vector(25 downto 0) := (others => 'X'); -- address
			avs_s0_read          : in  std_logic                     := 'X';             -- read
			avs_s0_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			avs_s0_write         : in  std_logic                     := 'X';             -- write
			avs_s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_s0_readdatavalid : out std_logic;                                        -- readdatavalid
			avs_s0_waitrequest   : out std_logic;                                        -- waitrequest
			avs_s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			avs_s0_burstcount    : in  std_logic_vector(6 downto 0)  := (others => 'X'); -- burstcount
			avm_m0_address       : out std_logic_vector(31 downto 0);                    -- address
			avm_m0_read          : out std_logic;                                        -- read
			avm_m0_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			avm_m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			avm_m0_write         : out std_logic;                                        -- write
			avm_m0_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			avm_m0_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			avm_m0_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			avm_m0_burstcount    : out std_logic_vector(6 downto 0);                     -- burstcount
			avs_cntl_address     : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- address
			avs_cntl_read        : in  std_logic                     := 'X';             -- read
			avs_cntl_readdata    : out std_logic_vector(63 downto 0);                    -- readdata
			avs_cntl_write       : in  std_logic                     := 'X';             -- write
			avs_cntl_writedata   : in  std_logic_vector(63 downto 0) := (others => 'X'); -- writedata
			avs_cntl_byteenable  : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- byteenable
		);
	end component altera_address_span_extender;

	component soc_system_hps_0 is
		generic (
			F2S_Width : integer := 2;
			S2F_Width : integer := 2
		);
		port (
			mem_a                    : out   std_logic_vector(14 downto 0);                    -- mem_a
			mem_ba                   : out   std_logic_vector(2 downto 0);                     -- mem_ba
			mem_ck                   : out   std_logic;                                        -- mem_ck
			mem_ck_n                 : out   std_logic;                                        -- mem_ck_n
			mem_cke                  : out   std_logic;                                        -- mem_cke
			mem_cs_n                 : out   std_logic;                                        -- mem_cs_n
			mem_ras_n                : out   std_logic;                                        -- mem_ras_n
			mem_cas_n                : out   std_logic;                                        -- mem_cas_n
			mem_we_n                 : out   std_logic;                                        -- mem_we_n
			mem_reset_n              : out   std_logic;                                        -- mem_reset_n
			mem_dq                   : inout std_logic_vector(31 downto 0) := (others => 'X'); -- mem_dq
			mem_dqs                  : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs
			mem_dqs_n                : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs_n
			mem_odt                  : out   std_logic;                                        -- mem_odt
			mem_dm                   : out   std_logic_vector(3 downto 0);                     -- mem_dm
			oct_rzqin                : in    std_logic                     := 'X';             -- oct_rzqin
			hps_io_emac1_inst_TX_CLK : out   std_logic;                                        -- hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0   : out   std_logic;                                        -- hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1   : out   std_logic;                                        -- hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2   : out   std_logic;                                        -- hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3   : out   std_logic;                                        -- hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO   : inout std_logic                     := 'X';             -- hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC    : out   std_logic;                                        -- hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL : out   std_logic;                                        -- hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD3
			hps_io_sdio_inst_CMD     : inout std_logic                     := 'X';             -- hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK     : out   std_logic;                                        -- hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D3
			hps_io_usb1_inst_D0      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D0
			hps_io_usb1_inst_D1      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D1
			hps_io_usb1_inst_D2      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D2
			hps_io_usb1_inst_D3      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D3
			hps_io_usb1_inst_D4      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D4
			hps_io_usb1_inst_D5      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D5
			hps_io_usb1_inst_D6      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D6
			hps_io_usb1_inst_D7      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D7
			hps_io_usb1_inst_CLK     : in    std_logic                     := 'X';             -- hps_io_usb1_inst_CLK
			hps_io_usb1_inst_STP     : out   std_logic;                                        -- hps_io_usb1_inst_STP
			hps_io_usb1_inst_DIR     : in    std_logic                     := 'X';             -- hps_io_usb1_inst_DIR
			hps_io_usb1_inst_NXT     : in    std_logic                     := 'X';             -- hps_io_usb1_inst_NXT
			hps_io_spim1_inst_CLK    : out   std_logic;                                        -- hps_io_spim1_inst_CLK
			hps_io_spim1_inst_MOSI   : out   std_logic;                                        -- hps_io_spim1_inst_MOSI
			hps_io_spim1_inst_MISO   : in    std_logic                     := 'X';             -- hps_io_spim1_inst_MISO
			hps_io_spim1_inst_SS0    : out   std_logic;                                        -- hps_io_spim1_inst_SS0
			hps_io_uart0_inst_RX     : in    std_logic                     := 'X';             -- hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     : out   std_logic;                                        -- hps_io_uart0_inst_TX
			hps_io_i2c0_inst_SDA     : inout std_logic                     := 'X';             -- hps_io_i2c0_inst_SDA
			hps_io_i2c0_inst_SCL     : inout std_logic                     := 'X';             -- hps_io_i2c0_inst_SCL
			hps_io_i2c1_inst_SDA     : inout std_logic                     := 'X';             -- hps_io_i2c1_inst_SDA
			hps_io_i2c1_inst_SCL     : inout std_logic                     := 'X';             -- hps_io_i2c1_inst_SCL
			hps_io_gpio_inst_GPIO09  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO09
			hps_io_gpio_inst_GPIO35  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO35
			hps_io_gpio_inst_GPIO40  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO40
			hps_io_gpio_inst_GPIO53  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO53
			hps_io_gpio_inst_GPIO54  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO54
			hps_io_gpio_inst_GPIO61  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO61
			h2f_rst_n                : out   std_logic;                                        -- reset_n
			f2h_sdram0_clk           : in    std_logic                     := 'X';             -- clk
			f2h_sdram0_ADDRESS       : in    std_logic_vector(29 downto 0) := (others => 'X'); -- address
			f2h_sdram0_BURSTCOUNT    : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- burstcount
			f2h_sdram0_WAITREQUEST   : out   std_logic;                                        -- waitrequest
			f2h_sdram0_READDATA      : out   std_logic_vector(31 downto 0);                    -- readdata
			f2h_sdram0_READDATAVALID : out   std_logic;                                        -- readdatavalid
			f2h_sdram0_READ          : in    std_logic                     := 'X';             -- read
			f2h_sdram0_WRITEDATA     : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			f2h_sdram0_BYTEENABLE    : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			f2h_sdram0_WRITE         : in    std_logic                     := 'X'              -- write
		);
	end component soc_system_hps_0;

	component soc_system_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component soc_system_jtag_uart_0;

	component soc_system_nios2_gen2_0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(30 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(30 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component soc_system_nios2_gen2_0;

	component soc_system_onchip_memory2_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component soc_system_onchip_memory2_0;

	component soc_system_pio_leds is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component soc_system_pio_leds;

	component soc_system_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                        : in  std_logic                     := 'X';             -- clk
			LCD_controller_0_reset_reset_bridge_in_reset_reset   : in  std_logic                     := 'X';             -- reset
			pio_leds_reset_reset_bridge_in_reset_reset           : in  std_logic                     := 'X';             -- reset
			LCD_controller_0_avalon_master_address               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			LCD_controller_0_avalon_master_waitrequest           : out std_logic;                                        -- waitrequest
			LCD_controller_0_avalon_master_burstcount            : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- burstcount
			LCD_controller_0_avalon_master_read                  : in  std_logic                     := 'X';             -- read
			LCD_controller_0_avalon_master_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			LCD_controller_0_avalon_master_readdatavalid         : out std_logic;                                        -- readdatavalid
			nios2_gen2_0_data_master_address                     : in  std_logic_vector(30 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_data_master_waitrequest                 : out std_logic;                                        -- waitrequest
			nios2_gen2_0_data_master_byteenable                  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_gen2_0_data_master_read                        : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_data_master_readdata                    : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_gen2_0_data_master_readdatavalid               : out std_logic;                                        -- readdatavalid
			nios2_gen2_0_data_master_write                       : in  std_logic                     := 'X';             -- write
			nios2_gen2_0_data_master_writedata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_gen2_0_data_master_debugaccess                 : in  std_logic                     := 'X';             -- debugaccess
			nios2_gen2_0_instruction_master_address              : in  std_logic_vector(30 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_instruction_master_waitrequest          : out std_logic;                                        -- waitrequest
			nios2_gen2_0_instruction_master_read                 : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_instruction_master_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_gen2_0_instruction_master_readdatavalid        : out std_logic;                                        -- readdatavalid
			address_span_extender_0_windowed_slave_address       : out std_logic_vector(25 downto 0);                    -- address
			address_span_extender_0_windowed_slave_write         : out std_logic;                                        -- write
			address_span_extender_0_windowed_slave_read          : out std_logic;                                        -- read
			address_span_extender_0_windowed_slave_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			address_span_extender_0_windowed_slave_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			address_span_extender_0_windowed_slave_burstcount    : out std_logic_vector(6 downto 0);                     -- burstcount
			address_span_extender_0_windowed_slave_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			address_span_extender_0_windowed_slave_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			address_span_extender_0_windowed_slave_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_address                : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write                  : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read                   : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata              : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest            : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect             : out std_logic;                                        -- chipselect
			LCD_controller_0_as_address                          : out std_logic_vector(3 downto 0);                     -- address
			LCD_controller_0_as_write                            : out std_logic;                                        -- write
			LCD_controller_0_as_read                             : out std_logic;                                        -- read
			LCD_controller_0_as_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			LCD_controller_0_as_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			LCD_controller_0_as_chipselect                       : out std_logic;                                        -- chipselect
			nios2_gen2_0_debug_mem_slave_address                 : out std_logic_vector(8 downto 0);                     -- address
			nios2_gen2_0_debug_mem_slave_write                   : out std_logic;                                        -- write
			nios2_gen2_0_debug_mem_slave_read                    : out std_logic;                                        -- read
			nios2_gen2_0_debug_mem_slave_readdata                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_gen2_0_debug_mem_slave_writedata               : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_gen2_0_debug_mem_slave_byteenable              : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest             : in  std_logic                     := 'X';             -- waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess             : out std_logic;                                        -- debugaccess
			onchip_memory2_0_s1_address                          : out std_logic_vector(14 downto 0);                    -- address
			onchip_memory2_0_s1_write                            : out std_logic;                                        -- write
			onchip_memory2_0_s1_readdata                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_memory2_0_s1_writedata                        : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_memory2_0_s1_byteenable                       : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_memory2_0_s1_chipselect                       : out std_logic;                                        -- chipselect
			onchip_memory2_0_s1_clken                            : out std_logic;                                        -- clken
			pio_leds_s1_address                                  : out std_logic_vector(1 downto 0);                     -- address
			pio_leds_s1_write                                    : out std_logic;                                        -- write
			pio_leds_s1_readdata                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_leds_s1_writedata                                : out std_logic_vector(31 downto 0);                    -- writedata
			pio_leds_s1_chipselect                               : out std_logic                                         -- chipselect
		);
	end component soc_system_mm_interconnect_0;

	component soc_system_mm_interconnect_1 is
		port (
			clk_0_clk_clk                                                      : in  std_logic                     := 'X';             -- clk
			address_span_extender_0_reset_reset_bridge_in_reset_reset          : in  std_logic                     := 'X';             -- reset
			hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			address_span_extender_0_expanded_master_address                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			address_span_extender_0_expanded_master_waitrequest                : out std_logic;                                        -- waitrequest
			address_span_extender_0_expanded_master_burstcount                 : in  std_logic_vector(6 downto 0)  := (others => 'X'); -- burstcount
			address_span_extender_0_expanded_master_byteenable                 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			address_span_extender_0_expanded_master_read                       : in  std_logic                     := 'X';             -- read
			address_span_extender_0_expanded_master_readdata                   : out std_logic_vector(31 downto 0);                    -- readdata
			address_span_extender_0_expanded_master_readdatavalid              : out std_logic;                                        -- readdatavalid
			address_span_extender_0_expanded_master_write                      : in  std_logic                     := 'X';             -- write
			address_span_extender_0_expanded_master_writedata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			hps_0_f2h_sdram0_data_address                                      : out std_logic_vector(29 downto 0);                    -- address
			hps_0_f2h_sdram0_data_write                                        : out std_logic;                                        -- write
			hps_0_f2h_sdram0_data_read                                         : out std_logic;                                        -- read
			hps_0_f2h_sdram0_data_readdata                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hps_0_f2h_sdram0_data_writedata                                    : out std_logic_vector(31 downto 0);                    -- writedata
			hps_0_f2h_sdram0_data_burstcount                                   : out std_logic_vector(7 downto 0);                     -- burstcount
			hps_0_f2h_sdram0_data_byteenable                                   : out std_logic_vector(3 downto 0);                     -- byteenable
			hps_0_f2h_sdram0_data_readdatavalid                                : in  std_logic                     := 'X';             -- readdatavalid
			hps_0_f2h_sdram0_data_waitrequest                                  : in  std_logic                     := 'X'              -- waitrequest
		);
	end component soc_system_mm_interconnect_1;

	component soc_system_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component soc_system_irq_mapper;

	component soc_system_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			reset_in2      : in  std_logic := 'X'; -- reset_in2.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component soc_system_rst_controller;

	component soc_system_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component soc_system_rst_controller_001;

	component soc_system_rst_controller_002 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component soc_system_rst_controller_002;

	signal lcd_controller_0_avalon_master_readdata                                : std_logic_vector(31 downto 0); -- mm_interconnect_0:LCD_controller_0_avalon_master_readdata -> LCD_controller_0:AM_readdata
	signal lcd_controller_0_avalon_master_waitrequest                             : std_logic;                     -- mm_interconnect_0:LCD_controller_0_avalon_master_waitrequest -> LCD_controller_0:AM_waitRQ
	signal lcd_controller_0_avalon_master_address                                 : std_logic_vector(31 downto 0); -- LCD_controller_0:AM_address -> mm_interconnect_0:LCD_controller_0_avalon_master_address
	signal lcd_controller_0_avalon_master_read                                    : std_logic;                     -- LCD_controller_0:AM_read -> mm_interconnect_0:LCD_controller_0_avalon_master_read
	signal lcd_controller_0_avalon_master_readdatavalid                           : std_logic;                     -- mm_interconnect_0:LCD_controller_0_avalon_master_readdatavalid -> LCD_controller_0:AM_Rddatavalid
	signal lcd_controller_0_avalon_master_burstcount                              : std_logic_vector(7 downto 0);  -- LCD_controller_0:AM_BurstCount -> mm_interconnect_0:LCD_controller_0_avalon_master_burstcount
	signal nios2_gen2_0_data_master_readdata                                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	signal nios2_gen2_0_data_master_waitrequest                                   : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	signal nios2_gen2_0_data_master_debugaccess                                   : std_logic;                     -- nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	signal nios2_gen2_0_data_master_address                                       : std_logic_vector(30 downto 0); -- nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	signal nios2_gen2_0_data_master_byteenable                                    : std_logic_vector(3 downto 0);  -- nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	signal nios2_gen2_0_data_master_read                                          : std_logic;                     -- nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	signal nios2_gen2_0_data_master_readdatavalid                                 : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_data_master_readdatavalid -> nios2_gen2_0:d_readdatavalid
	signal nios2_gen2_0_data_master_write                                         : std_logic;                     -- nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	signal nios2_gen2_0_data_master_writedata                                     : std_logic_vector(31 downto 0); -- nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	signal nios2_gen2_0_instruction_master_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	signal nios2_gen2_0_instruction_master_waitrequest                            : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	signal nios2_gen2_0_instruction_master_address                                : std_logic_vector(30 downto 0); -- nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	signal nios2_gen2_0_instruction_master_read                                   : std_logic;                     -- nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	signal nios2_gen2_0_instruction_master_readdatavalid                          : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_instruction_master_readdatavalid -> nios2_gen2_0:i_readdatavalid
	signal mm_interconnect_0_lcd_controller_0_as_chipselect                       : std_logic;                     -- mm_interconnect_0:LCD_controller_0_as_chipselect -> LCD_controller_0:AS_CS
	signal mm_interconnect_0_lcd_controller_0_as_readdata                         : std_logic_vector(31 downto 0); -- LCD_controller_0:AS_readdata -> mm_interconnect_0:LCD_controller_0_as_readdata
	signal mm_interconnect_0_lcd_controller_0_as_address                          : std_logic_vector(3 downto 0);  -- mm_interconnect_0:LCD_controller_0_as_address -> LCD_controller_0:AS_address
	signal mm_interconnect_0_lcd_controller_0_as_read                             : std_logic;                     -- mm_interconnect_0:LCD_controller_0_as_read -> LCD_controller_0:AS_read
	signal mm_interconnect_0_lcd_controller_0_as_write                            : std_logic;                     -- mm_interconnect_0:LCD_controller_0_as_write -> LCD_controller_0:AS_write
	signal mm_interconnect_0_lcd_controller_0_as_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:LCD_controller_0_as_writedata -> LCD_controller_0:AS_writedata
	signal mm_interconnect_0_pio_leds_s1_chipselect                               : std_logic;                     -- mm_interconnect_0:pio_leds_s1_chipselect -> pio_leds:chipselect
	signal mm_interconnect_0_pio_leds_s1_readdata                                 : std_logic_vector(31 downto 0); -- pio_leds:readdata -> mm_interconnect_0:pio_leds_s1_readdata
	signal mm_interconnect_0_pio_leds_s1_address                                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_leds_s1_address -> pio_leds:address
	signal mm_interconnect_0_pio_leds_s1_write                                    : std_logic;                     -- mm_interconnect_0:pio_leds_s1_write -> mm_interconnect_0_pio_leds_s1_write:in
	signal mm_interconnect_0_pio_leds_s1_writedata                                : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_leds_s1_writedata -> pio_leds:writedata
	signal mm_interconnect_0_address_span_extender_0_windowed_slave_readdata      : std_logic_vector(31 downto 0); -- address_span_extender_0:avs_s0_readdata -> mm_interconnect_0:address_span_extender_0_windowed_slave_readdata
	signal mm_interconnect_0_address_span_extender_0_windowed_slave_waitrequest   : std_logic;                     -- address_span_extender_0:avs_s0_waitrequest -> mm_interconnect_0:address_span_extender_0_windowed_slave_waitrequest
	signal mm_interconnect_0_address_span_extender_0_windowed_slave_address       : std_logic_vector(25 downto 0); -- mm_interconnect_0:address_span_extender_0_windowed_slave_address -> address_span_extender_0:avs_s0_address
	signal mm_interconnect_0_address_span_extender_0_windowed_slave_read          : std_logic;                     -- mm_interconnect_0:address_span_extender_0_windowed_slave_read -> address_span_extender_0:avs_s0_read
	signal mm_interconnect_0_address_span_extender_0_windowed_slave_byteenable    : std_logic_vector(3 downto 0);  -- mm_interconnect_0:address_span_extender_0_windowed_slave_byteenable -> address_span_extender_0:avs_s0_byteenable
	signal mm_interconnect_0_address_span_extender_0_windowed_slave_readdatavalid : std_logic;                     -- address_span_extender_0:avs_s0_readdatavalid -> mm_interconnect_0:address_span_extender_0_windowed_slave_readdatavalid
	signal mm_interconnect_0_address_span_extender_0_windowed_slave_write         : std_logic;                     -- mm_interconnect_0:address_span_extender_0_windowed_slave_write -> address_span_extender_0:avs_s0_write
	signal mm_interconnect_0_address_span_extender_0_windowed_slave_writedata     : std_logic_vector(31 downto 0); -- mm_interconnect_0:address_span_extender_0_windowed_slave_writedata -> address_span_extender_0:avs_s0_writedata
	signal mm_interconnect_0_address_span_extender_0_windowed_slave_burstcount    : std_logic_vector(6 downto 0);  -- mm_interconnect_0:address_span_extender_0_windowed_slave_burstcount -> address_span_extender_0:avs_s0_burstcount
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect             : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata               : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest            : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address                : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read                   : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write                  : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata              : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata                : std_logic_vector(31 downto 0); -- nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest             : std_logic;                     -- nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess             : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address                 : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read                    : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable              : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write                   : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata               : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	signal mm_interconnect_0_onchip_memory2_0_s1_readdata                         : std_logic_vector(31 downto 0); -- onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	signal mm_interconnect_0_onchip_memory2_0_s1_address                          : std_logic_vector(14 downto 0); -- mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	signal mm_interconnect_0_onchip_memory2_0_s1_byteenable                       : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	signal mm_interconnect_0_onchip_memory2_0_s1_write                            : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	signal mm_interconnect_0_onchip_memory2_0_s1_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	signal mm_interconnect_0_onchip_memory2_0_s1_clken                            : std_logic;                     -- mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	signal address_span_extender_0_expanded_master_waitrequest                    : std_logic;                     -- mm_interconnect_1:address_span_extender_0_expanded_master_waitrequest -> address_span_extender_0:avm_m0_waitrequest
	signal address_span_extender_0_expanded_master_readdata                       : std_logic_vector(31 downto 0); -- mm_interconnect_1:address_span_extender_0_expanded_master_readdata -> address_span_extender_0:avm_m0_readdata
	signal address_span_extender_0_expanded_master_address                        : std_logic_vector(31 downto 0); -- address_span_extender_0:avm_m0_address -> mm_interconnect_1:address_span_extender_0_expanded_master_address
	signal address_span_extender_0_expanded_master_read                           : std_logic;                     -- address_span_extender_0:avm_m0_read -> mm_interconnect_1:address_span_extender_0_expanded_master_read
	signal address_span_extender_0_expanded_master_byteenable                     : std_logic_vector(3 downto 0);  -- address_span_extender_0:avm_m0_byteenable -> mm_interconnect_1:address_span_extender_0_expanded_master_byteenable
	signal address_span_extender_0_expanded_master_readdatavalid                  : std_logic;                     -- mm_interconnect_1:address_span_extender_0_expanded_master_readdatavalid -> address_span_extender_0:avm_m0_readdatavalid
	signal address_span_extender_0_expanded_master_write                          : std_logic;                     -- address_span_extender_0:avm_m0_write -> mm_interconnect_1:address_span_extender_0_expanded_master_write
	signal address_span_extender_0_expanded_master_writedata                      : std_logic_vector(31 downto 0); -- address_span_extender_0:avm_m0_writedata -> mm_interconnect_1:address_span_extender_0_expanded_master_writedata
	signal address_span_extender_0_expanded_master_burstcount                     : std_logic_vector(6 downto 0);  -- address_span_extender_0:avm_m0_burstcount -> mm_interconnect_1:address_span_extender_0_expanded_master_burstcount
	signal mm_interconnect_1_hps_0_f2h_sdram0_data_readdata                       : std_logic_vector(31 downto 0); -- hps_0:f2h_sdram0_READDATA -> mm_interconnect_1:hps_0_f2h_sdram0_data_readdata
	signal mm_interconnect_1_hps_0_f2h_sdram0_data_waitrequest                    : std_logic;                     -- hps_0:f2h_sdram0_WAITREQUEST -> mm_interconnect_1:hps_0_f2h_sdram0_data_waitrequest
	signal mm_interconnect_1_hps_0_f2h_sdram0_data_address                        : std_logic_vector(29 downto 0); -- mm_interconnect_1:hps_0_f2h_sdram0_data_address -> hps_0:f2h_sdram0_ADDRESS
	signal mm_interconnect_1_hps_0_f2h_sdram0_data_read                           : std_logic;                     -- mm_interconnect_1:hps_0_f2h_sdram0_data_read -> hps_0:f2h_sdram0_READ
	signal mm_interconnect_1_hps_0_f2h_sdram0_data_byteenable                     : std_logic_vector(3 downto 0);  -- mm_interconnect_1:hps_0_f2h_sdram0_data_byteenable -> hps_0:f2h_sdram0_BYTEENABLE
	signal mm_interconnect_1_hps_0_f2h_sdram0_data_readdatavalid                  : std_logic;                     -- hps_0:f2h_sdram0_READDATAVALID -> mm_interconnect_1:hps_0_f2h_sdram0_data_readdatavalid
	signal mm_interconnect_1_hps_0_f2h_sdram0_data_write                          : std_logic;                     -- mm_interconnect_1:hps_0_f2h_sdram0_data_write -> hps_0:f2h_sdram0_WRITE
	signal mm_interconnect_1_hps_0_f2h_sdram0_data_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_1:hps_0_f2h_sdram0_data_writedata -> hps_0:f2h_sdram0_WRITEDATA
	signal mm_interconnect_1_hps_0_f2h_sdram0_data_burstcount                     : std_logic_vector(7 downto 0);  -- mm_interconnect_1:hps_0_f2h_sdram0_data_burstcount -> hps_0:f2h_sdram0_BURSTCOUNT
	signal irq_mapper_receiver0_irq                                               : std_logic;                     -- LCD_controller_0:AS_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                               : std_logic;                     -- jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	signal nios2_gen2_0_irq_irq                                                   : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_gen2_0:irq
	signal rst_controller_reset_out_reset                                         : std_logic;                     -- rst_controller:reset_out -> [address_span_extender_0:reset, irq_mapper:reset, mm_interconnect_0:LCD_controller_0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:address_span_extender_0_reset_reset_bridge_in_reset_reset, onchip_memory2_0:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                                     : std_logic;                     -- rst_controller:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	signal nios2_gen2_0_debug_reset_request_reset                                 : std_logic;                     -- nios2_gen2_0:debug_reset_request -> rst_controller:reset_in1
	signal hps_0_h2f_reset_reset                                                  : std_logic;                     -- hps_0:h2f_rst_n -> hps_0_h2f_reset_reset:in
	signal rst_controller_001_reset_out_reset                                     : std_logic;                     -- rst_controller_001:reset_out -> [mm_interconnect_0:pio_leds_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in]
	signal rst_controller_002_reset_out_reset                                     : std_logic;                     -- rst_controller_002:reset_out -> mm_interconnect_1:hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset_reset
	signal reset_reset_n_ports_inv                                                : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal mm_interconnect_0_pio_leds_s1_write_ports_inv                          : std_logic;                     -- mm_interconnect_0_pio_leds_s1_write:inv -> pio_leds:write_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv         : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv        : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal rst_controller_reset_out_reset_ports_inv                               : std_logic;                     -- rst_controller_reset_out_reset:inv -> [LCD_controller_0:nReset, jtag_uart_0:rst_n, nios2_gen2_0:reset_n]
	signal hps_0_h2f_reset_reset_ports_inv                                        : std_logic;                     -- hps_0_h2f_reset_reset:inv -> [rst_controller:reset_in2, rst_controller_001:reset_in1, rst_controller_002:reset_in0]
	signal rst_controller_001_reset_out_reset_ports_inv                           : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> pio_leds:reset_n

begin

	lcd_controller_0 : component LT24_controller
		port map (
			clk            => clk_clk,                                          --            clock.clk
			nReset         => rst_controller_reset_out_reset_ports_inv,         --            reset.reset_n
			AM_address     => lcd_controller_0_avalon_master_address,           --    avalon_master.address
			AM_read        => lcd_controller_0_avalon_master_read,              --                 .read
			AM_readdata    => lcd_controller_0_avalon_master_readdata,          --                 .readdata
			AM_waitRQ      => lcd_controller_0_avalon_master_waitrequest,       --                 .waitrequest
			AM_BurstCount  => lcd_controller_0_avalon_master_burstcount,        --                 .burstcount
			AM_Rddatavalid => lcd_controller_0_avalon_master_readdatavalid,     --                 .readdatavalid
			CS_N           => lcd_controller_0_conduit_end_export_cs_n,         --      conduit_end.export_cs_n
			DATA           => lcd_controller_0_conduit_end_export_data,         --                 .export_data
			D_C_N          => lcd_controller_0_conduit_end_export_d_c_n,        --                 .export_d_c_n
			LCD_ON         => lcd_controller_0_conduit_end_export_lcd_on,       --                 .export_lcd_on
			RD_N           => lcd_controller_0_conduit_end_export_rd_n,         --                 .export_rd_n
			RESET_N        => lcd_controller_0_conduit_end_export_reset_n,      --                 .export_reset_n
			WR_N           => lcd_controller_0_conduit_end_export_wr_n,         --                 .export_wr_n
			AS_address     => mm_interconnect_0_lcd_controller_0_as_address,    --               as.address
			AS_write       => mm_interconnect_0_lcd_controller_0_as_write,      --                 .write
			AS_writedata   => mm_interconnect_0_lcd_controller_0_as_writedata,  --                 .writedata
			AS_read        => mm_interconnect_0_lcd_controller_0_as_read,       --                 .read
			AS_readdata    => mm_interconnect_0_lcd_controller_0_as_readdata,   --                 .readdata
			AS_CS          => mm_interconnect_0_lcd_controller_0_as_chipselect, --                 .chipselect
			AS_irq         => irq_mapper_receiver0_irq                          -- interrupt_sender.irq
		);

	address_span_extender_0 : component altera_address_span_extender
		generic map (
			DATA_WIDTH           => 32,
			BYTEENABLE_WIDTH     => 4,
			MASTER_ADDRESS_WIDTH => 32,
			SLAVE_ADDRESS_WIDTH  => 26,
			SLAVE_ADDRESS_SHIFT  => 2,
			BURSTCOUNT_WIDTH     => 7,
			CNTL_ADDRESS_WIDTH   => 1,
			SUB_WINDOW_COUNT     => 1,
			MASTER_ADDRESS_DEF   => "0000000000000000000000000000000000110000000000000000000000000000"
		)
		port map (
			clk                  => clk_clk,                                                                --           clock.clk
			reset                => rst_controller_reset_out_reset,                                         --           reset.reset
			avs_s0_address       => mm_interconnect_0_address_span_extender_0_windowed_slave_address,       --  windowed_slave.address
			avs_s0_read          => mm_interconnect_0_address_span_extender_0_windowed_slave_read,          --                .read
			avs_s0_readdata      => mm_interconnect_0_address_span_extender_0_windowed_slave_readdata,      --                .readdata
			avs_s0_write         => mm_interconnect_0_address_span_extender_0_windowed_slave_write,         --                .write
			avs_s0_writedata     => mm_interconnect_0_address_span_extender_0_windowed_slave_writedata,     --                .writedata
			avs_s0_readdatavalid => mm_interconnect_0_address_span_extender_0_windowed_slave_readdatavalid, --                .readdatavalid
			avs_s0_waitrequest   => mm_interconnect_0_address_span_extender_0_windowed_slave_waitrequest,   --                .waitrequest
			avs_s0_byteenable    => mm_interconnect_0_address_span_extender_0_windowed_slave_byteenable,    --                .byteenable
			avs_s0_burstcount    => mm_interconnect_0_address_span_extender_0_windowed_slave_burstcount,    --                .burstcount
			avm_m0_address       => address_span_extender_0_expanded_master_address,                        -- expanded_master.address
			avm_m0_read          => address_span_extender_0_expanded_master_read,                           --                .read
			avm_m0_waitrequest   => address_span_extender_0_expanded_master_waitrequest,                    --                .waitrequest
			avm_m0_readdata      => address_span_extender_0_expanded_master_readdata,                       --                .readdata
			avm_m0_write         => address_span_extender_0_expanded_master_write,                          --                .write
			avm_m0_writedata     => address_span_extender_0_expanded_master_writedata,                      --                .writedata
			avm_m0_readdatavalid => address_span_extender_0_expanded_master_readdatavalid,                  --                .readdatavalid
			avm_m0_byteenable    => address_span_extender_0_expanded_master_byteenable,                     --                .byteenable
			avm_m0_burstcount    => address_span_extender_0_expanded_master_burstcount,                     --                .burstcount
			avs_cntl_address     => "0",                                                                    --     (terminated)
			avs_cntl_read        => '0',                                                                    --     (terminated)
			avs_cntl_readdata    => open,                                                                   --     (terminated)
			avs_cntl_write       => '0',                                                                    --     (terminated)
			avs_cntl_writedata   => "0000000000000000000000000000000000000000000000000000000000000000",     --     (terminated)
			avs_cntl_byteenable  => "00000000"                                                              --     (terminated)
		);

	hps_0 : component soc_system_hps_0
		generic map (
			F2S_Width => 0,
			S2F_Width => 0
		)
		port map (
			mem_a                    => hps_0_ddr_mem_a,                                       --           memory.mem_a
			mem_ba                   => hps_0_ddr_mem_ba,                                      --                 .mem_ba
			mem_ck                   => hps_0_ddr_mem_ck,                                      --                 .mem_ck
			mem_ck_n                 => hps_0_ddr_mem_ck_n,                                    --                 .mem_ck_n
			mem_cke                  => hps_0_ddr_mem_cke,                                     --                 .mem_cke
			mem_cs_n                 => hps_0_ddr_mem_cs_n,                                    --                 .mem_cs_n
			mem_ras_n                => hps_0_ddr_mem_ras_n,                                   --                 .mem_ras_n
			mem_cas_n                => hps_0_ddr_mem_cas_n,                                   --                 .mem_cas_n
			mem_we_n                 => hps_0_ddr_mem_we_n,                                    --                 .mem_we_n
			mem_reset_n              => hps_0_ddr_mem_reset_n,                                 --                 .mem_reset_n
			mem_dq                   => hps_0_ddr_mem_dq,                                      --                 .mem_dq
			mem_dqs                  => hps_0_ddr_mem_dqs,                                     --                 .mem_dqs
			mem_dqs_n                => hps_0_ddr_mem_dqs_n,                                   --                 .mem_dqs_n
			mem_odt                  => hps_0_ddr_mem_odt,                                     --                 .mem_odt
			mem_dm                   => hps_0_ddr_mem_dm,                                      --                 .mem_dm
			oct_rzqin                => hps_0_ddr_oct_rzqin,                                   --                 .oct_rzqin
			hps_io_emac1_inst_TX_CLK => hps_0_io_hps_io_emac1_inst_TX_CLK,                     --           hps_io.hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0   => hps_0_io_hps_io_emac1_inst_TXD0,                       --                 .hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1   => hps_0_io_hps_io_emac1_inst_TXD1,                       --                 .hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2   => hps_0_io_hps_io_emac1_inst_TXD2,                       --                 .hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3   => hps_0_io_hps_io_emac1_inst_TXD3,                       --                 .hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0   => hps_0_io_hps_io_emac1_inst_RXD0,                       --                 .hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO   => hps_0_io_hps_io_emac1_inst_MDIO,                       --                 .hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC    => hps_0_io_hps_io_emac1_inst_MDC,                        --                 .hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL => hps_0_io_hps_io_emac1_inst_RX_CTL,                     --                 .hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL => hps_0_io_hps_io_emac1_inst_TX_CTL,                     --                 .hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK => hps_0_io_hps_io_emac1_inst_RX_CLK,                     --                 .hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1   => hps_0_io_hps_io_emac1_inst_RXD1,                       --                 .hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2   => hps_0_io_hps_io_emac1_inst_RXD2,                       --                 .hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3   => hps_0_io_hps_io_emac1_inst_RXD3,                       --                 .hps_io_emac1_inst_RXD3
			hps_io_sdio_inst_CMD     => hps_0_io_hps_io_sdio_inst_CMD,                         --                 .hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0      => hps_0_io_hps_io_sdio_inst_D0,                          --                 .hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1      => hps_0_io_hps_io_sdio_inst_D1,                          --                 .hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK     => hps_0_io_hps_io_sdio_inst_CLK,                         --                 .hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2      => hps_0_io_hps_io_sdio_inst_D2,                          --                 .hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3      => hps_0_io_hps_io_sdio_inst_D3,                          --                 .hps_io_sdio_inst_D3
			hps_io_usb1_inst_D0      => hps_0_io_hps_io_usb1_inst_D0,                          --                 .hps_io_usb1_inst_D0
			hps_io_usb1_inst_D1      => hps_0_io_hps_io_usb1_inst_D1,                          --                 .hps_io_usb1_inst_D1
			hps_io_usb1_inst_D2      => hps_0_io_hps_io_usb1_inst_D2,                          --                 .hps_io_usb1_inst_D2
			hps_io_usb1_inst_D3      => hps_0_io_hps_io_usb1_inst_D3,                          --                 .hps_io_usb1_inst_D3
			hps_io_usb1_inst_D4      => hps_0_io_hps_io_usb1_inst_D4,                          --                 .hps_io_usb1_inst_D4
			hps_io_usb1_inst_D5      => hps_0_io_hps_io_usb1_inst_D5,                          --                 .hps_io_usb1_inst_D5
			hps_io_usb1_inst_D6      => hps_0_io_hps_io_usb1_inst_D6,                          --                 .hps_io_usb1_inst_D6
			hps_io_usb1_inst_D7      => hps_0_io_hps_io_usb1_inst_D7,                          --                 .hps_io_usb1_inst_D7
			hps_io_usb1_inst_CLK     => hps_0_io_hps_io_usb1_inst_CLK,                         --                 .hps_io_usb1_inst_CLK
			hps_io_usb1_inst_STP     => hps_0_io_hps_io_usb1_inst_STP,                         --                 .hps_io_usb1_inst_STP
			hps_io_usb1_inst_DIR     => hps_0_io_hps_io_usb1_inst_DIR,                         --                 .hps_io_usb1_inst_DIR
			hps_io_usb1_inst_NXT     => hps_0_io_hps_io_usb1_inst_NXT,                         --                 .hps_io_usb1_inst_NXT
			hps_io_spim1_inst_CLK    => hps_0_io_hps_io_spim1_inst_CLK,                        --                 .hps_io_spim1_inst_CLK
			hps_io_spim1_inst_MOSI   => hps_0_io_hps_io_spim1_inst_MOSI,                       --                 .hps_io_spim1_inst_MOSI
			hps_io_spim1_inst_MISO   => hps_0_io_hps_io_spim1_inst_MISO,                       --                 .hps_io_spim1_inst_MISO
			hps_io_spim1_inst_SS0    => hps_0_io_hps_io_spim1_inst_SS0,                        --                 .hps_io_spim1_inst_SS0
			hps_io_uart0_inst_RX     => hps_0_io_hps_io_uart0_inst_RX,                         --                 .hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     => hps_0_io_hps_io_uart0_inst_TX,                         --                 .hps_io_uart0_inst_TX
			hps_io_i2c0_inst_SDA     => hps_0_io_hps_io_i2c0_inst_SDA,                         --                 .hps_io_i2c0_inst_SDA
			hps_io_i2c0_inst_SCL     => hps_0_io_hps_io_i2c0_inst_SCL,                         --                 .hps_io_i2c0_inst_SCL
			hps_io_i2c1_inst_SDA     => hps_0_io_hps_io_i2c1_inst_SDA,                         --                 .hps_io_i2c1_inst_SDA
			hps_io_i2c1_inst_SCL     => hps_0_io_hps_io_i2c1_inst_SCL,                         --                 .hps_io_i2c1_inst_SCL
			hps_io_gpio_inst_GPIO09  => hps_0_io_hps_io_gpio_inst_GPIO09,                      --                 .hps_io_gpio_inst_GPIO09
			hps_io_gpio_inst_GPIO35  => hps_0_io_hps_io_gpio_inst_GPIO35,                      --                 .hps_io_gpio_inst_GPIO35
			hps_io_gpio_inst_GPIO40  => hps_0_io_hps_io_gpio_inst_GPIO40,                      --                 .hps_io_gpio_inst_GPIO40
			hps_io_gpio_inst_GPIO53  => hps_0_io_hps_io_gpio_inst_GPIO53,                      --                 .hps_io_gpio_inst_GPIO53
			hps_io_gpio_inst_GPIO54  => hps_0_io_hps_io_gpio_inst_GPIO54,                      --                 .hps_io_gpio_inst_GPIO54
			hps_io_gpio_inst_GPIO61  => hps_0_io_hps_io_gpio_inst_GPIO61,                      --                 .hps_io_gpio_inst_GPIO61
			h2f_rst_n                => hps_0_h2f_reset_reset,                                 --        h2f_reset.reset_n
			f2h_sdram0_clk           => clk_clk,                                               -- f2h_sdram0_clock.clk
			f2h_sdram0_ADDRESS       => mm_interconnect_1_hps_0_f2h_sdram0_data_address,       --  f2h_sdram0_data.address
			f2h_sdram0_BURSTCOUNT    => mm_interconnect_1_hps_0_f2h_sdram0_data_burstcount,    --                 .burstcount
			f2h_sdram0_WAITREQUEST   => mm_interconnect_1_hps_0_f2h_sdram0_data_waitrequest,   --                 .waitrequest
			f2h_sdram0_READDATA      => mm_interconnect_1_hps_0_f2h_sdram0_data_readdata,      --                 .readdata
			f2h_sdram0_READDATAVALID => mm_interconnect_1_hps_0_f2h_sdram0_data_readdatavalid, --                 .readdatavalid
			f2h_sdram0_READ          => mm_interconnect_1_hps_0_f2h_sdram0_data_read,          --                 .read
			f2h_sdram0_WRITEDATA     => mm_interconnect_1_hps_0_f2h_sdram0_data_writedata,     --                 .writedata
			f2h_sdram0_BYTEENABLE    => mm_interconnect_1_hps_0_f2h_sdram0_data_byteenable,    --                 .byteenable
			f2h_sdram0_WRITE         => mm_interconnect_1_hps_0_f2h_sdram0_data_write          --                 .write
		);

	jtag_uart_0 : component soc_system_jtag_uart_0
		port map (
			clk            => clk_clk,                                                         --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                        --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver1_irq                                         --               irq.irq
		);

	nios2_gen2_0 : component soc_system_nios2_gen2_0
		port map (
			clk                                 => clk_clk,                                                    --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,                   --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                         --                          .reset_req
			d_address                           => nios2_gen2_0_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_gen2_0_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_gen2_0_data_master_read,                              --                          .read
			d_readdata                          => nios2_gen2_0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_gen2_0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_gen2_0_data_master_write,                             --                          .write
			d_writedata                         => nios2_gen2_0_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => nios2_gen2_0_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => nios2_gen2_0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_gen2_0_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_gen2_0_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_gen2_0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_gen2_0_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => nios2_gen2_0_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => nios2_gen2_0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2_gen2_0_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                        -- custom_instruction_master.readra
		);

	onchip_memory2_0 : component soc_system_onchip_memory2_0
		port map (
			clk        => clk_clk,                                          --   clk1.clk
			address    => mm_interconnect_0_onchip_memory2_0_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_memory2_0_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_memory2_0_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_memory2_0_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_memory2_0_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_memory2_0_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_memory2_0_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                   -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,               --       .reset_req
			freeze     => '0'                                               -- (terminated)
		);

	pio_leds : component soc_system_pio_leds
		port map (
			clk        => clk_clk,                                       --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_pio_leds_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_leds_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_leds_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_leds_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_leds_s1_readdata,        --                    .readdata
			out_port   => pio_leds_external_connection_export            -- external_connection.export
		);

	mm_interconnect_0 : component soc_system_mm_interconnect_0
		port map (
			clk_0_clk_clk                                        => clk_clk,                                                                --                                    clk_0_clk.clk
			LCD_controller_0_reset_reset_bridge_in_reset_reset   => rst_controller_reset_out_reset,                                         -- LCD_controller_0_reset_reset_bridge_in_reset.reset
			pio_leds_reset_reset_bridge_in_reset_reset           => rst_controller_001_reset_out_reset,                                     --         pio_leds_reset_reset_bridge_in_reset.reset
			LCD_controller_0_avalon_master_address               => lcd_controller_0_avalon_master_address,                                 --               LCD_controller_0_avalon_master.address
			LCD_controller_0_avalon_master_waitrequest           => lcd_controller_0_avalon_master_waitrequest,                             --                                             .waitrequest
			LCD_controller_0_avalon_master_burstcount            => lcd_controller_0_avalon_master_burstcount,                              --                                             .burstcount
			LCD_controller_0_avalon_master_read                  => lcd_controller_0_avalon_master_read,                                    --                                             .read
			LCD_controller_0_avalon_master_readdata              => lcd_controller_0_avalon_master_readdata,                                --                                             .readdata
			LCD_controller_0_avalon_master_readdatavalid         => lcd_controller_0_avalon_master_readdatavalid,                           --                                             .readdatavalid
			nios2_gen2_0_data_master_address                     => nios2_gen2_0_data_master_address,                                       --                     nios2_gen2_0_data_master.address
			nios2_gen2_0_data_master_waitrequest                 => nios2_gen2_0_data_master_waitrequest,                                   --                                             .waitrequest
			nios2_gen2_0_data_master_byteenable                  => nios2_gen2_0_data_master_byteenable,                                    --                                             .byteenable
			nios2_gen2_0_data_master_read                        => nios2_gen2_0_data_master_read,                                          --                                             .read
			nios2_gen2_0_data_master_readdata                    => nios2_gen2_0_data_master_readdata,                                      --                                             .readdata
			nios2_gen2_0_data_master_readdatavalid               => nios2_gen2_0_data_master_readdatavalid,                                 --                                             .readdatavalid
			nios2_gen2_0_data_master_write                       => nios2_gen2_0_data_master_write,                                         --                                             .write
			nios2_gen2_0_data_master_writedata                   => nios2_gen2_0_data_master_writedata,                                     --                                             .writedata
			nios2_gen2_0_data_master_debugaccess                 => nios2_gen2_0_data_master_debugaccess,                                   --                                             .debugaccess
			nios2_gen2_0_instruction_master_address              => nios2_gen2_0_instruction_master_address,                                --              nios2_gen2_0_instruction_master.address
			nios2_gen2_0_instruction_master_waitrequest          => nios2_gen2_0_instruction_master_waitrequest,                            --                                             .waitrequest
			nios2_gen2_0_instruction_master_read                 => nios2_gen2_0_instruction_master_read,                                   --                                             .read
			nios2_gen2_0_instruction_master_readdata             => nios2_gen2_0_instruction_master_readdata,                               --                                             .readdata
			nios2_gen2_0_instruction_master_readdatavalid        => nios2_gen2_0_instruction_master_readdatavalid,                          --                                             .readdatavalid
			address_span_extender_0_windowed_slave_address       => mm_interconnect_0_address_span_extender_0_windowed_slave_address,       --       address_span_extender_0_windowed_slave.address
			address_span_extender_0_windowed_slave_write         => mm_interconnect_0_address_span_extender_0_windowed_slave_write,         --                                             .write
			address_span_extender_0_windowed_slave_read          => mm_interconnect_0_address_span_extender_0_windowed_slave_read,          --                                             .read
			address_span_extender_0_windowed_slave_readdata      => mm_interconnect_0_address_span_extender_0_windowed_slave_readdata,      --                                             .readdata
			address_span_extender_0_windowed_slave_writedata     => mm_interconnect_0_address_span_extender_0_windowed_slave_writedata,     --                                             .writedata
			address_span_extender_0_windowed_slave_burstcount    => mm_interconnect_0_address_span_extender_0_windowed_slave_burstcount,    --                                             .burstcount
			address_span_extender_0_windowed_slave_byteenable    => mm_interconnect_0_address_span_extender_0_windowed_slave_byteenable,    --                                             .byteenable
			address_span_extender_0_windowed_slave_readdatavalid => mm_interconnect_0_address_span_extender_0_windowed_slave_readdatavalid, --                                             .readdatavalid
			address_span_extender_0_windowed_slave_waitrequest   => mm_interconnect_0_address_span_extender_0_windowed_slave_waitrequest,   --                                             .waitrequest
			jtag_uart_0_avalon_jtag_slave_address                => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address,                --                jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write                  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write,                  --                                             .write
			jtag_uart_0_avalon_jtag_slave_read                   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read,                   --                                             .read
			jtag_uart_0_avalon_jtag_slave_readdata               => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,               --                                             .readdata
			jtag_uart_0_avalon_jtag_slave_writedata              => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,              --                                             .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest            => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,            --                                             .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect             => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,             --                                             .chipselect
			LCD_controller_0_as_address                          => mm_interconnect_0_lcd_controller_0_as_address,                          --                          LCD_controller_0_as.address
			LCD_controller_0_as_write                            => mm_interconnect_0_lcd_controller_0_as_write,                            --                                             .write
			LCD_controller_0_as_read                             => mm_interconnect_0_lcd_controller_0_as_read,                             --                                             .read
			LCD_controller_0_as_readdata                         => mm_interconnect_0_lcd_controller_0_as_readdata,                         --                                             .readdata
			LCD_controller_0_as_writedata                        => mm_interconnect_0_lcd_controller_0_as_writedata,                        --                                             .writedata
			LCD_controller_0_as_chipselect                       => mm_interconnect_0_lcd_controller_0_as_chipselect,                       --                                             .chipselect
			nios2_gen2_0_debug_mem_slave_address                 => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,                 --                 nios2_gen2_0_debug_mem_slave.address
			nios2_gen2_0_debug_mem_slave_write                   => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,                   --                                             .write
			nios2_gen2_0_debug_mem_slave_read                    => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,                    --                                             .read
			nios2_gen2_0_debug_mem_slave_readdata                => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,                --                                             .readdata
			nios2_gen2_0_debug_mem_slave_writedata               => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,               --                                             .writedata
			nios2_gen2_0_debug_mem_slave_byteenable              => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,              --                                             .byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest,             --                                             .waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess,             --                                             .debugaccess
			onchip_memory2_0_s1_address                          => mm_interconnect_0_onchip_memory2_0_s1_address,                          --                          onchip_memory2_0_s1.address
			onchip_memory2_0_s1_write                            => mm_interconnect_0_onchip_memory2_0_s1_write,                            --                                             .write
			onchip_memory2_0_s1_readdata                         => mm_interconnect_0_onchip_memory2_0_s1_readdata,                         --                                             .readdata
			onchip_memory2_0_s1_writedata                        => mm_interconnect_0_onchip_memory2_0_s1_writedata,                        --                                             .writedata
			onchip_memory2_0_s1_byteenable                       => mm_interconnect_0_onchip_memory2_0_s1_byteenable,                       --                                             .byteenable
			onchip_memory2_0_s1_chipselect                       => mm_interconnect_0_onchip_memory2_0_s1_chipselect,                       --                                             .chipselect
			onchip_memory2_0_s1_clken                            => mm_interconnect_0_onchip_memory2_0_s1_clken,                            --                                             .clken
			pio_leds_s1_address                                  => mm_interconnect_0_pio_leds_s1_address,                                  --                                  pio_leds_s1.address
			pio_leds_s1_write                                    => mm_interconnect_0_pio_leds_s1_write,                                    --                                             .write
			pio_leds_s1_readdata                                 => mm_interconnect_0_pio_leds_s1_readdata,                                 --                                             .readdata
			pio_leds_s1_writedata                                => mm_interconnect_0_pio_leds_s1_writedata,                                --                                             .writedata
			pio_leds_s1_chipselect                               => mm_interconnect_0_pio_leds_s1_chipselect                                --                                             .chipselect
		);

	mm_interconnect_1 : component soc_system_mm_interconnect_1
		port map (
			clk_0_clk_clk                                                      => clk_clk,                                               --                                                    clk_0_clk.clk
			address_span_extender_0_reset_reset_bridge_in_reset_reset          => rst_controller_reset_out_reset,                        --          address_span_extender_0_reset_reset_bridge_in_reset.reset
			hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset_reset => rst_controller_002_reset_out_reset,                    -- hps_0_f2h_sdram0_data_translator_reset_reset_bridge_in_reset.reset
			address_span_extender_0_expanded_master_address                    => address_span_extender_0_expanded_master_address,       --                      address_span_extender_0_expanded_master.address
			address_span_extender_0_expanded_master_waitrequest                => address_span_extender_0_expanded_master_waitrequest,   --                                                             .waitrequest
			address_span_extender_0_expanded_master_burstcount                 => address_span_extender_0_expanded_master_burstcount,    --                                                             .burstcount
			address_span_extender_0_expanded_master_byteenable                 => address_span_extender_0_expanded_master_byteenable,    --                                                             .byteenable
			address_span_extender_0_expanded_master_read                       => address_span_extender_0_expanded_master_read,          --                                                             .read
			address_span_extender_0_expanded_master_readdata                   => address_span_extender_0_expanded_master_readdata,      --                                                             .readdata
			address_span_extender_0_expanded_master_readdatavalid              => address_span_extender_0_expanded_master_readdatavalid, --                                                             .readdatavalid
			address_span_extender_0_expanded_master_write                      => address_span_extender_0_expanded_master_write,         --                                                             .write
			address_span_extender_0_expanded_master_writedata                  => address_span_extender_0_expanded_master_writedata,     --                                                             .writedata
			hps_0_f2h_sdram0_data_address                                      => mm_interconnect_1_hps_0_f2h_sdram0_data_address,       --                                        hps_0_f2h_sdram0_data.address
			hps_0_f2h_sdram0_data_write                                        => mm_interconnect_1_hps_0_f2h_sdram0_data_write,         --                                                             .write
			hps_0_f2h_sdram0_data_read                                         => mm_interconnect_1_hps_0_f2h_sdram0_data_read,          --                                                             .read
			hps_0_f2h_sdram0_data_readdata                                     => mm_interconnect_1_hps_0_f2h_sdram0_data_readdata,      --                                                             .readdata
			hps_0_f2h_sdram0_data_writedata                                    => mm_interconnect_1_hps_0_f2h_sdram0_data_writedata,     --                                                             .writedata
			hps_0_f2h_sdram0_data_burstcount                                   => mm_interconnect_1_hps_0_f2h_sdram0_data_burstcount,    --                                                             .burstcount
			hps_0_f2h_sdram0_data_byteenable                                   => mm_interconnect_1_hps_0_f2h_sdram0_data_byteenable,    --                                                             .byteenable
			hps_0_f2h_sdram0_data_readdatavalid                                => mm_interconnect_1_hps_0_f2h_sdram0_data_readdatavalid, --                                                             .readdatavalid
			hps_0_f2h_sdram0_data_waitrequest                                  => mm_interconnect_1_hps_0_f2h_sdram0_data_waitrequest    --                                                             .waitrequest
		);

	irq_mapper : component soc_system_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			sender_irq    => nios2_gen2_0_irq_irq            --    sender.irq
		);

	rst_controller : component soc_system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 3,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			reset_in1      => nios2_gen2_0_debug_reset_request_reset, -- reset_in1.reset
			reset_in2      => hps_0_h2f_reset_reset_ports_inv,        -- reset_in2.reset
			clk            => clk_clk,                                --       clk.clk
			reset_out      => rst_controller_reset_out_reset,         -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,     --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_001 : component soc_system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => hps_0_h2f_reset_reset_ports_inv,    -- reset_in1.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_002 : component soc_system_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => hps_0_h2f_reset_reset_ports_inv,    -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_pio_leds_s1_write_ports_inv <= not mm_interconnect_0_pio_leds_s1_write;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	hps_0_h2f_reset_reset_ports_inv <= not hps_0_h2f_reset_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of soc_system
