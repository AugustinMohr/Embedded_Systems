library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity Segment_7 is

	port(
	
		clk		: in std_logic;
		nReset	: in std_logic;
		
		
		--Internal interface (i.e. Avalon slave).
		
		--External interface (i.e. conduit)
		
	);
end Segment_7;

architecture comp of Segment_7 is


signal 



begin

	
end comp;	
					