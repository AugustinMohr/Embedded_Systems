
module unsaved (
	clk_clk,
	reset_reset_n,
	enable_writeresponsevalid_n);	

	input		clk_clk;
	input		reset_reset_n;
	output		enable_writeresponsevalid_n;
endmodule
