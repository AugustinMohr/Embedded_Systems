library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity Avalon_Master is

	port(
	
		clk		: in std_logic;
		nReset	: in std_logic;
		
		
		--Internal interface (i.e. Avalon slave).
		
		--External interface (i.e. conduit)
		
	);
end Avalon_Master;

architecture comp of Avalon_Master is


signal 



begin

	
end comp;	
					