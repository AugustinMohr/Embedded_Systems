
module system2_1 (
	clk_clk,
	custom_pio_0_external_connection_export,
	reset_reset_n);	

	input		clk_clk;
	inout	[7:0]	custom_pio_0_external_connection_export;
	input		reset_reset_n;
endmodule
